// pruebaS7.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module pruebaS7 (
		input  wire [1:0] btn_pin_export,     //     btn_pin.export
		input  wire       clk_clk,            //         clk.clk
		output wire [7:0] led_pin_export,     //     led_pin.export
		input  wire       reset_reset_n,      //       reset.reset_n
		output wire [6:0] seg_7_0_pin_export, // seg_7_0_pin.export
		output wire [6:0] seg_7_1_pin_export, // seg_7_1_pin.export
		output wire [6:0] seg_7_2_pin_export, // seg_7_2_pin.export
		output wire [6:0] seg_7_3_pin_export, // seg_7_3_pin.export
		output wire [6:0] seg_7_4_pin_export, // seg_7_4_pin.export
		input  wire [7:0] sw_pin_export       //      sw_pin.export
	);

	wire  [31:0] nios_cpu_data_master_readdata;                          // mm_interconnect_0:NIOS_CPU_data_master_readdata -> NIOS_CPU:d_readdata
	wire         nios_cpu_data_master_waitrequest;                       // mm_interconnect_0:NIOS_CPU_data_master_waitrequest -> NIOS_CPU:d_waitrequest
	wire         nios_cpu_data_master_debugaccess;                       // NIOS_CPU:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:NIOS_CPU_data_master_debugaccess
	wire  [13:0] nios_cpu_data_master_address;                           // NIOS_CPU:d_address -> mm_interconnect_0:NIOS_CPU_data_master_address
	wire   [3:0] nios_cpu_data_master_byteenable;                        // NIOS_CPU:d_byteenable -> mm_interconnect_0:NIOS_CPU_data_master_byteenable
	wire         nios_cpu_data_master_read;                              // NIOS_CPU:d_read -> mm_interconnect_0:NIOS_CPU_data_master_read
	wire         nios_cpu_data_master_write;                             // NIOS_CPU:d_write -> mm_interconnect_0:NIOS_CPU_data_master_write
	wire  [31:0] nios_cpu_data_master_writedata;                         // NIOS_CPU:d_writedata -> mm_interconnect_0:NIOS_CPU_data_master_writedata
	wire  [31:0] nios_cpu_instruction_master_readdata;                   // mm_interconnect_0:NIOS_CPU_instruction_master_readdata -> NIOS_CPU:i_readdata
	wire         nios_cpu_instruction_master_waitrequest;                // mm_interconnect_0:NIOS_CPU_instruction_master_waitrequest -> NIOS_CPU:i_waitrequest
	wire  [13:0] nios_cpu_instruction_master_address;                    // NIOS_CPU:i_address -> mm_interconnect_0:NIOS_CPU_instruction_master_address
	wire         nios_cpu_instruction_master_read;                       // NIOS_CPU:i_read -> mm_interconnect_0:NIOS_CPU_instruction_master_read
	wire         mm_interconnect_0_uart_avalon_jtag_slave_chipselect;    // mm_interconnect_0:UART_avalon_jtag_slave_chipselect -> UART:av_chipselect
	wire  [31:0] mm_interconnect_0_uart_avalon_jtag_slave_readdata;      // UART:av_readdata -> mm_interconnect_0:UART_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_uart_avalon_jtag_slave_waitrequest;   // UART:av_waitrequest -> mm_interconnect_0:UART_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_uart_avalon_jtag_slave_address;       // mm_interconnect_0:UART_avalon_jtag_slave_address -> UART:av_address
	wire         mm_interconnect_0_uart_avalon_jtag_slave_read;          // mm_interconnect_0:UART_avalon_jtag_slave_read -> UART:av_read_n
	wire         mm_interconnect_0_uart_avalon_jtag_slave_write;         // mm_interconnect_0:UART_avalon_jtag_slave_write -> UART:av_write_n
	wire  [31:0] mm_interconnect_0_uart_avalon_jtag_slave_writedata;     // mm_interconnect_0:UART_avalon_jtag_slave_writedata -> UART:av_writedata
	wire  [31:0] mm_interconnect_0_nios_cpu_debug_mem_slave_readdata;    // NIOS_CPU:debug_mem_slave_readdata -> mm_interconnect_0:NIOS_CPU_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios_cpu_debug_mem_slave_waitrequest; // NIOS_CPU:debug_mem_slave_waitrequest -> mm_interconnect_0:NIOS_CPU_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios_cpu_debug_mem_slave_debugaccess; // mm_interconnect_0:NIOS_CPU_debug_mem_slave_debugaccess -> NIOS_CPU:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios_cpu_debug_mem_slave_address;     // mm_interconnect_0:NIOS_CPU_debug_mem_slave_address -> NIOS_CPU:debug_mem_slave_address
	wire         mm_interconnect_0_nios_cpu_debug_mem_slave_read;        // mm_interconnect_0:NIOS_CPU_debug_mem_slave_read -> NIOS_CPU:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios_cpu_debug_mem_slave_byteenable;  // mm_interconnect_0:NIOS_CPU_debug_mem_slave_byteenable -> NIOS_CPU:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios_cpu_debug_mem_slave_write;       // mm_interconnect_0:NIOS_CPU_debug_mem_slave_write -> NIOS_CPU:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios_cpu_debug_mem_slave_writedata;   // mm_interconnect_0:NIOS_CPU_debug_mem_slave_writedata -> NIOS_CPU:debug_mem_slave_writedata
	wire         mm_interconnect_0_ram_s1_chipselect;                    // mm_interconnect_0:RAM_s1_chipselect -> RAM:chipselect
	wire  [31:0] mm_interconnect_0_ram_s1_readdata;                      // RAM:readdata -> mm_interconnect_0:RAM_s1_readdata
	wire   [9:0] mm_interconnect_0_ram_s1_address;                       // mm_interconnect_0:RAM_s1_address -> RAM:address
	wire   [3:0] mm_interconnect_0_ram_s1_byteenable;                    // mm_interconnect_0:RAM_s1_byteenable -> RAM:byteenable
	wire         mm_interconnect_0_ram_s1_write;                         // mm_interconnect_0:RAM_s1_write -> RAM:write
	wire  [31:0] mm_interconnect_0_ram_s1_writedata;                     // mm_interconnect_0:RAM_s1_writedata -> RAM:writedata
	wire         mm_interconnect_0_ram_s1_clken;                         // mm_interconnect_0:RAM_s1_clken -> RAM:clken
	wire         mm_interconnect_0_led_s1_chipselect;                    // mm_interconnect_0:LED_s1_chipselect -> LED:chipselect
	wire  [31:0] mm_interconnect_0_led_s1_readdata;                      // LED:readdata -> mm_interconnect_0:LED_s1_readdata
	wire   [1:0] mm_interconnect_0_led_s1_address;                       // mm_interconnect_0:LED_s1_address -> LED:address
	wire         mm_interconnect_0_led_s1_write;                         // mm_interconnect_0:LED_s1_write -> LED:write_n
	wire  [31:0] mm_interconnect_0_led_s1_writedata;                     // mm_interconnect_0:LED_s1_writedata -> LED:writedata
	wire  [31:0] mm_interconnect_0_sw_s1_readdata;                       // SW:readdata -> mm_interconnect_0:SW_s1_readdata
	wire   [1:0] mm_interconnect_0_sw_s1_address;                        // mm_interconnect_0:SW_s1_address -> SW:address
	wire  [31:0] mm_interconnect_0_btn_s1_readdata;                      // BTN:readdata -> mm_interconnect_0:BTN_s1_readdata
	wire   [1:0] mm_interconnect_0_btn_s1_address;                       // mm_interconnect_0:BTN_s1_address -> BTN:address
	wire         mm_interconnect_0_seg_7_0_s1_chipselect;                // mm_interconnect_0:SEG_7_0_s1_chipselect -> SEG_7_0:chipselect
	wire  [31:0] mm_interconnect_0_seg_7_0_s1_readdata;                  // SEG_7_0:readdata -> mm_interconnect_0:SEG_7_0_s1_readdata
	wire   [1:0] mm_interconnect_0_seg_7_0_s1_address;                   // mm_interconnect_0:SEG_7_0_s1_address -> SEG_7_0:address
	wire         mm_interconnect_0_seg_7_0_s1_write;                     // mm_interconnect_0:SEG_7_0_s1_write -> SEG_7_0:write_n
	wire  [31:0] mm_interconnect_0_seg_7_0_s1_writedata;                 // mm_interconnect_0:SEG_7_0_s1_writedata -> SEG_7_0:writedata
	wire         mm_interconnect_0_seg_7_1_s1_chipselect;                // mm_interconnect_0:SEG_7_1_s1_chipselect -> SEG_7_1:chipselect
	wire  [31:0] mm_interconnect_0_seg_7_1_s1_readdata;                  // SEG_7_1:readdata -> mm_interconnect_0:SEG_7_1_s1_readdata
	wire   [1:0] mm_interconnect_0_seg_7_1_s1_address;                   // mm_interconnect_0:SEG_7_1_s1_address -> SEG_7_1:address
	wire         mm_interconnect_0_seg_7_1_s1_write;                     // mm_interconnect_0:SEG_7_1_s1_write -> SEG_7_1:write_n
	wire  [31:0] mm_interconnect_0_seg_7_1_s1_writedata;                 // mm_interconnect_0:SEG_7_1_s1_writedata -> SEG_7_1:writedata
	wire         mm_interconnect_0_seg_7_2_s1_chipselect;                // mm_interconnect_0:SEG_7_2_s1_chipselect -> SEG_7_2:chipselect
	wire  [31:0] mm_interconnect_0_seg_7_2_s1_readdata;                  // SEG_7_2:readdata -> mm_interconnect_0:SEG_7_2_s1_readdata
	wire   [1:0] mm_interconnect_0_seg_7_2_s1_address;                   // mm_interconnect_0:SEG_7_2_s1_address -> SEG_7_2:address
	wire         mm_interconnect_0_seg_7_2_s1_write;                     // mm_interconnect_0:SEG_7_2_s1_write -> SEG_7_2:write_n
	wire  [31:0] mm_interconnect_0_seg_7_2_s1_writedata;                 // mm_interconnect_0:SEG_7_2_s1_writedata -> SEG_7_2:writedata
	wire         mm_interconnect_0_seg_7_3_s1_chipselect;                // mm_interconnect_0:SEG_7_3_s1_chipselect -> SEG_7_3:chipselect
	wire  [31:0] mm_interconnect_0_seg_7_3_s1_readdata;                  // SEG_7_3:readdata -> mm_interconnect_0:SEG_7_3_s1_readdata
	wire   [1:0] mm_interconnect_0_seg_7_3_s1_address;                   // mm_interconnect_0:SEG_7_3_s1_address -> SEG_7_3:address
	wire         mm_interconnect_0_seg_7_3_s1_write;                     // mm_interconnect_0:SEG_7_3_s1_write -> SEG_7_3:write_n
	wire  [31:0] mm_interconnect_0_seg_7_3_s1_writedata;                 // mm_interconnect_0:SEG_7_3_s1_writedata -> SEG_7_3:writedata
	wire         mm_interconnect_0_seg_7_4_s1_chipselect;                // mm_interconnect_0:SEG_7_4_s1_chipselect -> SEG_7_4:chipselect
	wire  [31:0] mm_interconnect_0_seg_7_4_s1_readdata;                  // SEG_7_4:readdata -> mm_interconnect_0:SEG_7_4_s1_readdata
	wire   [1:0] mm_interconnect_0_seg_7_4_s1_address;                   // mm_interconnect_0:SEG_7_4_s1_address -> SEG_7_4:address
	wire         mm_interconnect_0_seg_7_4_s1_write;                     // mm_interconnect_0:SEG_7_4_s1_write -> SEG_7_4:write_n
	wire  [31:0] mm_interconnect_0_seg_7_4_s1_writedata;                 // mm_interconnect_0:SEG_7_4_s1_writedata -> SEG_7_4:writedata
	wire         irq_mapper_receiver0_irq;                               // UART:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] nios_cpu_irq_irq;                                       // irq_mapper:sender_irq -> NIOS_CPU:irq
	wire         rst_controller_reset_out_reset;                         // rst_controller:reset_out -> [BTN:reset_n, LED:reset_n, NIOS_CPU:reset_n, RAM:reset, SEG_7_0:reset_n, SEG_7_1:reset_n, SEG_7_2:reset_n, SEG_7_3:reset_n, SEG_7_4:reset_n, SW:reset_n, UART:rst_n, irq_mapper:reset, mm_interconnect_0:NIOS_CPU_reset_reset_bridge_in_reset_reset, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                     // rst_controller:reset_req -> [NIOS_CPU:reset_req, RAM:reset_req, rst_translator:reset_req_in]

	pruebaS7_BTN btn (
		.clk      (clk_clk),                           //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),   //               reset.reset_n
		.address  (mm_interconnect_0_btn_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_btn_s1_readdata), //                    .readdata
		.in_port  (btn_pin_export)                     // external_connection.export
	);

	pruebaS7_LED led (
		.clk        (clk_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led_s1_readdata),   //                    .readdata
		.out_port   (led_pin_export)                       // external_connection.export
	);

	pruebaS7_NIOS_CPU nios_cpu (
		.clk                                 (clk_clk),                                                //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                        //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                     //                          .reset_req
		.d_address                           (nios_cpu_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios_cpu_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios_cpu_data_master_read),                              //                          .read
		.d_readdata                          (nios_cpu_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios_cpu_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios_cpu_data_master_write),                             //                          .write
		.d_writedata                         (nios_cpu_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios_cpu_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios_cpu_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios_cpu_instruction_master_read),                       //                          .read
		.i_readdata                          (nios_cpu_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios_cpu_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios_cpu_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                       //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios_cpu_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios_cpu_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios_cpu_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios_cpu_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios_cpu_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios_cpu_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios_cpu_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios_cpu_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                        // custom_instruction_master.readra
	);

	pruebaS7_RAM ram (
		.clk        (clk_clk),                             //   clk1.clk
		.address    (mm_interconnect_0_ram_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_ram_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_ram_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_ram_s1_write),      //       .write
		.readdata   (mm_interconnect_0_ram_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_ram_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_ram_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),      // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),  //       .reset_req
		.freeze     (1'b0)                                 // (terminated)
	);

	pruebaS7_SEG_7_0 seg_7_0 (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_seg_7_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_seg_7_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_seg_7_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_seg_7_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_seg_7_0_s1_readdata),   //                    .readdata
		.out_port   (seg_7_0_pin_export)                       // external_connection.export
	);

	pruebaS7_SEG_7_0 seg_7_1 (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_seg_7_1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_seg_7_1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_seg_7_1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_seg_7_1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_seg_7_1_s1_readdata),   //                    .readdata
		.out_port   (seg_7_1_pin_export)                       // external_connection.export
	);

	pruebaS7_SEG_7_0 seg_7_2 (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_seg_7_2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_seg_7_2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_seg_7_2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_seg_7_2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_seg_7_2_s1_readdata),   //                    .readdata
		.out_port   (seg_7_2_pin_export)                       // external_connection.export
	);

	pruebaS7_SEG_7_0 seg_7_3 (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_seg_7_3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_seg_7_3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_seg_7_3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_seg_7_3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_seg_7_3_s1_readdata),   //                    .readdata
		.out_port   (seg_7_3_pin_export)                       // external_connection.export
	);

	pruebaS7_SEG_7_0 seg_7_4 (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_seg_7_4_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_seg_7_4_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_seg_7_4_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_seg_7_4_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_seg_7_4_s1_readdata),   //                    .readdata
		.out_port   (seg_7_4_pin_export)                       // external_connection.export
	);

	pruebaS7_SW sw (
		.clk      (clk_clk),                          //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),  //               reset.reset_n
		.address  (mm_interconnect_0_sw_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_sw_s1_readdata), //                    .readdata
		.in_port  (sw_pin_export)                     // external_connection.export
	);

	pruebaS7_UART uart (
		.clk            (clk_clk),                                              //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                      //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                              //               irq.irq
	);

	pruebaS7_mm_interconnect_0 mm_interconnect_0 (
		.CLK_clk_clk                                (clk_clk),                                                //                              CLK_clk.clk
		.NIOS_CPU_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                         // NIOS_CPU_reset_reset_bridge_in_reset.reset
		.NIOS_CPU_data_master_address               (nios_cpu_data_master_address),                           //                 NIOS_CPU_data_master.address
		.NIOS_CPU_data_master_waitrequest           (nios_cpu_data_master_waitrequest),                       //                                     .waitrequest
		.NIOS_CPU_data_master_byteenable            (nios_cpu_data_master_byteenable),                        //                                     .byteenable
		.NIOS_CPU_data_master_read                  (nios_cpu_data_master_read),                              //                                     .read
		.NIOS_CPU_data_master_readdata              (nios_cpu_data_master_readdata),                          //                                     .readdata
		.NIOS_CPU_data_master_write                 (nios_cpu_data_master_write),                             //                                     .write
		.NIOS_CPU_data_master_writedata             (nios_cpu_data_master_writedata),                         //                                     .writedata
		.NIOS_CPU_data_master_debugaccess           (nios_cpu_data_master_debugaccess),                       //                                     .debugaccess
		.NIOS_CPU_instruction_master_address        (nios_cpu_instruction_master_address),                    //          NIOS_CPU_instruction_master.address
		.NIOS_CPU_instruction_master_waitrequest    (nios_cpu_instruction_master_waitrequest),                //                                     .waitrequest
		.NIOS_CPU_instruction_master_read           (nios_cpu_instruction_master_read),                       //                                     .read
		.NIOS_CPU_instruction_master_readdata       (nios_cpu_instruction_master_readdata),                   //                                     .readdata
		.BTN_s1_address                             (mm_interconnect_0_btn_s1_address),                       //                               BTN_s1.address
		.BTN_s1_readdata                            (mm_interconnect_0_btn_s1_readdata),                      //                                     .readdata
		.LED_s1_address                             (mm_interconnect_0_led_s1_address),                       //                               LED_s1.address
		.LED_s1_write                               (mm_interconnect_0_led_s1_write),                         //                                     .write
		.LED_s1_readdata                            (mm_interconnect_0_led_s1_readdata),                      //                                     .readdata
		.LED_s1_writedata                           (mm_interconnect_0_led_s1_writedata),                     //                                     .writedata
		.LED_s1_chipselect                          (mm_interconnect_0_led_s1_chipselect),                    //                                     .chipselect
		.NIOS_CPU_debug_mem_slave_address           (mm_interconnect_0_nios_cpu_debug_mem_slave_address),     //             NIOS_CPU_debug_mem_slave.address
		.NIOS_CPU_debug_mem_slave_write             (mm_interconnect_0_nios_cpu_debug_mem_slave_write),       //                                     .write
		.NIOS_CPU_debug_mem_slave_read              (mm_interconnect_0_nios_cpu_debug_mem_slave_read),        //                                     .read
		.NIOS_CPU_debug_mem_slave_readdata          (mm_interconnect_0_nios_cpu_debug_mem_slave_readdata),    //                                     .readdata
		.NIOS_CPU_debug_mem_slave_writedata         (mm_interconnect_0_nios_cpu_debug_mem_slave_writedata),   //                                     .writedata
		.NIOS_CPU_debug_mem_slave_byteenable        (mm_interconnect_0_nios_cpu_debug_mem_slave_byteenable),  //                                     .byteenable
		.NIOS_CPU_debug_mem_slave_waitrequest       (mm_interconnect_0_nios_cpu_debug_mem_slave_waitrequest), //                                     .waitrequest
		.NIOS_CPU_debug_mem_slave_debugaccess       (mm_interconnect_0_nios_cpu_debug_mem_slave_debugaccess), //                                     .debugaccess
		.RAM_s1_address                             (mm_interconnect_0_ram_s1_address),                       //                               RAM_s1.address
		.RAM_s1_write                               (mm_interconnect_0_ram_s1_write),                         //                                     .write
		.RAM_s1_readdata                            (mm_interconnect_0_ram_s1_readdata),                      //                                     .readdata
		.RAM_s1_writedata                           (mm_interconnect_0_ram_s1_writedata),                     //                                     .writedata
		.RAM_s1_byteenable                          (mm_interconnect_0_ram_s1_byteenable),                    //                                     .byteenable
		.RAM_s1_chipselect                          (mm_interconnect_0_ram_s1_chipselect),                    //                                     .chipselect
		.RAM_s1_clken                               (mm_interconnect_0_ram_s1_clken),                         //                                     .clken
		.SEG_7_0_s1_address                         (mm_interconnect_0_seg_7_0_s1_address),                   //                           SEG_7_0_s1.address
		.SEG_7_0_s1_write                           (mm_interconnect_0_seg_7_0_s1_write),                     //                                     .write
		.SEG_7_0_s1_readdata                        (mm_interconnect_0_seg_7_0_s1_readdata),                  //                                     .readdata
		.SEG_7_0_s1_writedata                       (mm_interconnect_0_seg_7_0_s1_writedata),                 //                                     .writedata
		.SEG_7_0_s1_chipselect                      (mm_interconnect_0_seg_7_0_s1_chipselect),                //                                     .chipselect
		.SEG_7_1_s1_address                         (mm_interconnect_0_seg_7_1_s1_address),                   //                           SEG_7_1_s1.address
		.SEG_7_1_s1_write                           (mm_interconnect_0_seg_7_1_s1_write),                     //                                     .write
		.SEG_7_1_s1_readdata                        (mm_interconnect_0_seg_7_1_s1_readdata),                  //                                     .readdata
		.SEG_7_1_s1_writedata                       (mm_interconnect_0_seg_7_1_s1_writedata),                 //                                     .writedata
		.SEG_7_1_s1_chipselect                      (mm_interconnect_0_seg_7_1_s1_chipselect),                //                                     .chipselect
		.SEG_7_2_s1_address                         (mm_interconnect_0_seg_7_2_s1_address),                   //                           SEG_7_2_s1.address
		.SEG_7_2_s1_write                           (mm_interconnect_0_seg_7_2_s1_write),                     //                                     .write
		.SEG_7_2_s1_readdata                        (mm_interconnect_0_seg_7_2_s1_readdata),                  //                                     .readdata
		.SEG_7_2_s1_writedata                       (mm_interconnect_0_seg_7_2_s1_writedata),                 //                                     .writedata
		.SEG_7_2_s1_chipselect                      (mm_interconnect_0_seg_7_2_s1_chipselect),                //                                     .chipselect
		.SEG_7_3_s1_address                         (mm_interconnect_0_seg_7_3_s1_address),                   //                           SEG_7_3_s1.address
		.SEG_7_3_s1_write                           (mm_interconnect_0_seg_7_3_s1_write),                     //                                     .write
		.SEG_7_3_s1_readdata                        (mm_interconnect_0_seg_7_3_s1_readdata),                  //                                     .readdata
		.SEG_7_3_s1_writedata                       (mm_interconnect_0_seg_7_3_s1_writedata),                 //                                     .writedata
		.SEG_7_3_s1_chipselect                      (mm_interconnect_0_seg_7_3_s1_chipselect),                //                                     .chipselect
		.SEG_7_4_s1_address                         (mm_interconnect_0_seg_7_4_s1_address),                   //                           SEG_7_4_s1.address
		.SEG_7_4_s1_write                           (mm_interconnect_0_seg_7_4_s1_write),                     //                                     .write
		.SEG_7_4_s1_readdata                        (mm_interconnect_0_seg_7_4_s1_readdata),                  //                                     .readdata
		.SEG_7_4_s1_writedata                       (mm_interconnect_0_seg_7_4_s1_writedata),                 //                                     .writedata
		.SEG_7_4_s1_chipselect                      (mm_interconnect_0_seg_7_4_s1_chipselect),                //                                     .chipselect
		.SW_s1_address                              (mm_interconnect_0_sw_s1_address),                        //                                SW_s1.address
		.SW_s1_readdata                             (mm_interconnect_0_sw_s1_readdata),                       //                                     .readdata
		.UART_avalon_jtag_slave_address             (mm_interconnect_0_uart_avalon_jtag_slave_address),       //               UART_avalon_jtag_slave.address
		.UART_avalon_jtag_slave_write               (mm_interconnect_0_uart_avalon_jtag_slave_write),         //                                     .write
		.UART_avalon_jtag_slave_read                (mm_interconnect_0_uart_avalon_jtag_slave_read),          //                                     .read
		.UART_avalon_jtag_slave_readdata            (mm_interconnect_0_uart_avalon_jtag_slave_readdata),      //                                     .readdata
		.UART_avalon_jtag_slave_writedata           (mm_interconnect_0_uart_avalon_jtag_slave_writedata),     //                                     .writedata
		.UART_avalon_jtag_slave_waitrequest         (mm_interconnect_0_uart_avalon_jtag_slave_waitrequest),   //                                     .waitrequest
		.UART_avalon_jtag_slave_chipselect          (mm_interconnect_0_uart_avalon_jtag_slave_chipselect)     //                                     .chipselect
	);

	pruebaS7_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (nios_cpu_irq_irq)                //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
